module add_significands (
    sig1_cc, sig2_a, co, sum
);

input [26:0] sig1_cc, sig2_a;
output logic co;
output logic [26:0] sum;

endmodule