/*
 * File: \normalize.sv
 * Project: c:\Users\Chuck\ECE571\final_project\RISC-V-Floating-Point-Processor\src\design\chuck_test_code
 * Created Date: Thursday, May 6th 2021, 11:36:37 pm
 * Author: Chuck Faber
 * -----
 * Last Modified: Mon May 10 2021
 * Modified By: Chuck Faber
 * -----
 * Copyright (c) 2021 Portland State University
 * 
 * Takes in the summed significands, and carry out from the ALU checks 
 * if normalization is necessary and performs the normalization shift necessary.
 * 
 * Outputs the normalized signficand, and the shift value (negative for
 * left shift, positive for right shift) which will be added to the exponent.
 * 
 * -----
 * HISTORY:
 * Date      	By	Comments
 * ----------	---	----------------------------------------------------------
 */

module normalize (
    sig, carryout, sig_norm, shift
);

input [23:0] sig;
input carryout;
output logic [23:0] sig_norm;
output logic [7:0] shift;

if (carryout) begin                     // If there is a carryout we need to shift just 1 to the right, and increment the exponent.
    sig_norm = sig >> 1;
    shift = 1;
end else begin                          // Else keep shifting to the left and decrementing exponent until there is a 1 in the MSB.
    shift = 0;
    while (sig[23] != 1'b1) begin
        sig = sig << 1;
        shift -= 1;
    end
    sig_norm = sig;
end

endmodule