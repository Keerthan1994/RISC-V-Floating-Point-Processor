import addpkg::*;

module top();
    initial begin
        FpUnpackTest(0.25);
        FpUnpackTest(100);

    end

endmodule